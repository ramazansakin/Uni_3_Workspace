`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 	    Mehmet Akif TAŞOVA
// 
// Create Date:    20:22:29 11/17/2013 
// Design Name: 
// Module Name:    ALU-32Bit 
// Project Name:   32 Bit ALU
// Target Devices: 
// Tool versions: 
// Description: 
//			
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module ALU32Bit();


endmodule
